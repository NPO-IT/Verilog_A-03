module Astra (
	input clk80,
	input clk100
);

endmodule
